module mux_8x1(out, i0, i1, i2, i3, i4, i5, i6, i7, s0, s1, s2);
output out; 
input i0, i1, i2, i3, i4, i5, i6, i7, s0, s1, s2;

assign out = (s2 == 0) ? ((s1 == 0) ? ((s0 == 0) ? i0 : i1) : ((s0 == 0) ? i2 : i3)) : ((s1 == 0) ? ((s0 == 0) ? i4 : i5) : ((s0 == 0) ? i6 : i7)); 
endmodule
