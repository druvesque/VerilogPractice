module tb;
     reg clk;
     initial begin
         clk = 0;
         forever #10 clk = ~clk;
     end

     initial begin
         #200;
         $finish;
     end
endmodule
