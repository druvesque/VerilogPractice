module tb;

reg i0, i1, i2, i3, i4, i5, i6, i7, s0, s1, s2;
wire out;
mux_8x1 m1(out, i0, i1, i2, i3, i4, i5, i6, i7, s0, s1, s2);

initial begin
i0 = 1; i1 = 0; i2 = 0; i3 = 0; i4 = 0; i5 = 0; i6 = 0; i7 = 0; s2 = 0; s1 = 0; s0 = 0;
#10;
i0 = 0; i1 = 1; i2 = 0; i3 = 0; i4 = 0; i5 = 0; i6 = 0; i7 = 0; s2 = 0; s1 = 0; s0 = 1;
#10;
i0 = 0; i1 = 0; i2 = 1; i3 = 0; i4 = 0; i5 = 0; i6 = 0; i7 = 0; s2 = 0; s1 = 1; s0 = 0;
#10
i0 = 0; i1 = 0; i2 = 0; i3 = 1; i4 = 0; i5 = 0; i6 = 0; i7 = 0; s2 = 0; s1 = 1; s0 = 1;
#10
i0 = 0; i1 = 0; i2 = 0; i3 = 0; i4 = 1; i5 = 0; i6 = 0; i7 = 0; s2 = 1; s1 = 0; s0 = 0;
#10;
i0 = 0; i1 = 0; i2 = 0; i3 = 0; i4 = 0; i5 = 1; i6 = 0; i7 = 0; s2 = 1; s1 = 0; s0 = 1;
#10;
i0 = 0; i1 = 0; i2 = 0; i3 = 0; i4 = 0; i5 = 0; i6 = 1; i7 = 0; s2 = 1; s1 = 1; s0 = 0;
#10;
i0 = 0; i1 = 0; i2 = 0; i3 = 0; i4 = 0; i5 = 0; i6 = 0; i7 = 1; s2 = 1; s1 = 1; s0 = 1; 

end

initial begin
$monitor("Time: %t, i0: %d, i1: %d, i2: %d, i3: %d, i4: %d, i5: %d, i6: %d, i7: %d, s0: %d, s1: %d, s0: %d, Output: %d", $time, i0, i1, i2, i3, i4, i5, i6, i7, s0, s1, s2, out);
end

initial begin
$dumpfile("mux.vcd");
$dumpvars(0, tb);
end

initial begin
#200;
$finish;
end

endmodule
