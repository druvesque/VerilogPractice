module or_gate(o, a, b);
    input a, b;
    output o;

    assign o = a | b;
endmodule
