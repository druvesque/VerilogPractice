module display(
    input clk,
    output reg [6:0] y
);
    integer count = 0;

    always @(posedge clk)
    begin
        count <= count + 1;
        $display("\n Count: %d", count);
    end

    always @(posedge clk) begin
        case (count)
            0: y <= 7'b0000001; 
            1: y <= 7'b1001111;
            2: y <= 7'b0010010;
            3: y <= 7'b0000110;
            4: y <= 7'b1001100;
            5: y <= 7'b0100100;
            6: y <= 7'b0100000;
            7: y <= 7'b0001111;
            8: y <= 7'b0000000;
            9: y <= 7'b0000100;
        endcase
    end
endmodule

module tb;
    reg clk = 0;
    wire [6:0] y;
    display d1(.clk(clk), .y(y));

    initial 
        forever #5 clk = ~clk;
    initial begin
        $monitor("Time: %g, Output: %b", $time, y);

        $dumpfile("wv.vcd");
        $dumpvars(0, tb);

        #200;
        $finish;
    end
endmodule
