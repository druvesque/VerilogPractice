module checksum(a, b);
    input [63:0] a;
    input [7:0] b;
    assign b=doChecksum(a);

    function [7:0] doCheckSum;
        input [63:0] DataArray;
        reg [15:0] temp1, temp2;
        begin
            temp1 = DataArray[15:0] ^ DataArray[31:16];
            temp2 = DataArray[63:48] ^ DataArray[47:32];
            doCheckSum = temp1[7:0] + temp2[7:0] ^ temp1[15:8] + temp2[15:8];
        end
    endfunction
endmodule

module checksum_tb;
    reg [63:0] a;
    reg [7:0] b;

endmodule
